module SieveOfEratosthenesTest ();

	logic clock, reset_n, done;
	logic [100:0] is_prime;

//	SieveOfEratosthenes dut(.*);

//	initial begin
//		clock = 0;
//		forever #5 clock = ~clock;
//	end

//	initial 
//	begin 
//		$dumpfile("SieveOfEratosthenesBaseline_tb.vcd");
//		$dumpvars(1,dut);
//		$dumpon;
//		reset_n = 0;
//		reset_n <= 1;
//		$display("%b",done);
//		while(done !== 1)
//		begin
//			@(posedge clock);
//		end
//		foreach(is_prime[j]) begin
//			if(!is_prime[j]) 
//			begin
//				$display("%d\n",j);
//			end
//		// end
//		$dumpoff;
//		#10 $finish;
	//end

endmodule